

-- THIS FILE WAS AUTOMATICALLY GENERERATED. DO NOT MODIY BY HAND
-- GENERERATED BY ... 
-- Date

--------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.numeric_std.all;
use std.env.all;


entity test_iir_TB is
end test_iir_TB;

architecture TB of test_iir_TB is

component test_iir is
port (
  DATA_IN : signed(15 downto 0);
  DATA_IN_VAL : std_logic;
  CLK : in std_logic;
  SRST : in std_logic;
  DATA_OUT : out signed(17 downto 0);
  DATA_OUT_VAL : out std_logic
);
end component;


signal CLK : std_logic := '0';
constant CLK_PERIOD : time := 10.0 ns;

signal DATA_IN : signed(15 downto 0);
signal DATA_IN_VAL : std_logic := '0';
signal DATA_OUT_VAL : std_logic;
signal DATA_OUT : signed(17 downto 0);
signal SRST : std_logic := '0';


type DATA_IN_ARRAY_T is array (natural range <>) of signed(15 downto 0);

constant DATA_IN_ARRAY : DATA_IN_ARRAY_T(0 to 899) :=
(0 => to_signed(32767, 16),
 1 => to_signed(32767, 16),
 2 => to_signed(32767, 16),
 3 => to_signed(32767, 16),
 4 => to_signed(32767, 16),
 5 => to_signed(32767, 16),
 6 => to_signed(32767, 16),
 7 => to_signed(32767, 16),
 8 => to_signed(32767, 16),
 9 => to_signed(32767, 16),
 10 => to_signed(32767, 16),
 11 => to_signed(32767, 16),
 12 => to_signed(32767, 16),
 13 => to_signed(32767, 16),
 14 => to_signed(32767, 16),
 15 => to_signed(32767, 16),
 16 => to_signed(32767, 16),
 17 => to_signed(32767, 16),
 18 => to_signed(32767, 16),
 19 => to_signed(32767, 16),
 20 => to_signed(32767, 16),
 21 => to_signed(32767, 16),
 22 => to_signed(32767, 16),
 23 => to_signed(32767, 16),
 24 => to_signed(32767, 16),
 25 => to_signed(32767, 16),
 26 => to_signed(32767, 16),
 27 => to_signed(32767, 16),
 28 => to_signed(32767, 16),
 29 => to_signed(32767, 16),
 30 => to_signed(32767, 16),
 31 => to_signed(32767, 16),
 32 => to_signed(32767, 16),
 33 => to_signed(32767, 16),
 34 => to_signed(32767, 16),
 35 => to_signed(32767, 16),
 36 => to_signed(32767, 16),
 37 => to_signed(32767, 16),
 38 => to_signed(32767, 16),
 39 => to_signed(32767, 16),
 40 => to_signed(32767, 16),
 41 => to_signed(32767, 16),
 42 => to_signed(32767, 16),
 43 => to_signed(32767, 16),
 44 => to_signed(32767, 16),
 45 => to_signed(32767, 16),
 46 => to_signed(32767, 16),
 47 => to_signed(32767, 16),
 48 => to_signed(32767, 16),
 49 => to_signed(32767, 16),
 50 => to_signed(32767, 16),
 51 => to_signed(32767, 16),
 52 => to_signed(32767, 16),
 53 => to_signed(32767, 16),
 54 => to_signed(32767, 16),
 55 => to_signed(32767, 16),
 56 => to_signed(32767, 16),
 57 => to_signed(32767, 16),
 58 => to_signed(32767, 16),
 59 => to_signed(32767, 16),
 60 => to_signed(32767, 16),
 61 => to_signed(32767, 16),
 62 => to_signed(32767, 16),
 63 => to_signed(32767, 16),
 64 => to_signed(32767, 16),
 65 => to_signed(32767, 16),
 66 => to_signed(32767, 16),
 67 => to_signed(32767, 16),
 68 => to_signed(32767, 16),
 69 => to_signed(32767, 16),
 70 => to_signed(32767, 16),
 71 => to_signed(32767, 16),
 72 => to_signed(32767, 16),
 73 => to_signed(32767, 16),
 74 => to_signed(32767, 16),
 75 => to_signed(32767, 16),
 76 => to_signed(32767, 16),
 77 => to_signed(32767, 16),
 78 => to_signed(32767, 16),
 79 => to_signed(32767, 16),
 80 => to_signed(32767, 16),
 81 => to_signed(32767, 16),
 82 => to_signed(32767, 16),
 83 => to_signed(32767, 16),
 84 => to_signed(32767, 16),
 85 => to_signed(32767, 16),
 86 => to_signed(32767, 16),
 87 => to_signed(32767, 16),
 88 => to_signed(32767, 16),
 89 => to_signed(32767, 16),
 90 => to_signed(32767, 16),
 91 => to_signed(32767, 16),
 92 => to_signed(32767, 16),
 93 => to_signed(32767, 16),
 94 => to_signed(32767, 16),
 95 => to_signed(32767, 16),
 96 => to_signed(32767, 16),
 97 => to_signed(32767, 16),
 98 => to_signed(32767, 16),
 99 => to_signed(32767, 16),
 100 => to_signed(32767, 16),
 101 => to_signed(32767, 16),
 102 => to_signed(32767, 16),
 103 => to_signed(32767, 16),
 104 => to_signed(32767, 16),
 105 => to_signed(32767, 16),
 106 => to_signed(32767, 16),
 107 => to_signed(32767, 16),
 108 => to_signed(32767, 16),
 109 => to_signed(32767, 16),
 110 => to_signed(32767, 16),
 111 => to_signed(32767, 16),
 112 => to_signed(32767, 16),
 113 => to_signed(32767, 16),
 114 => to_signed(32767, 16),
 115 => to_signed(32767, 16),
 116 => to_signed(32767, 16),
 117 => to_signed(32767, 16),
 118 => to_signed(32767, 16),
 119 => to_signed(32767, 16),
 120 => to_signed(32767, 16),
 121 => to_signed(32767, 16),
 122 => to_signed(32767, 16),
 123 => to_signed(32767, 16),
 124 => to_signed(32767, 16),
 125 => to_signed(32767, 16),
 126 => to_signed(32767, 16),
 127 => to_signed(32767, 16),
 128 => to_signed(32767, 16),
 129 => to_signed(32767, 16),
 130 => to_signed(32767, 16),
 131 => to_signed(32767, 16),
 132 => to_signed(32767, 16),
 133 => to_signed(32767, 16),
 134 => to_signed(32767, 16),
 135 => to_signed(32767, 16),
 136 => to_signed(32767, 16),
 137 => to_signed(32767, 16),
 138 => to_signed(32767, 16),
 139 => to_signed(32767, 16),
 140 => to_signed(32767, 16),
 141 => to_signed(32767, 16),
 142 => to_signed(32767, 16),
 143 => to_signed(32767, 16),
 144 => to_signed(32767, 16),
 145 => to_signed(32767, 16),
 146 => to_signed(32767, 16),
 147 => to_signed(32767, 16),
 148 => to_signed(32767, 16),
 149 => to_signed(32767, 16),
 150 => to_signed(32767, 16),
 151 => to_signed(32767, 16),
 152 => to_signed(32767, 16),
 153 => to_signed(32767, 16),
 154 => to_signed(32767, 16),
 155 => to_signed(32767, 16),
 156 => to_signed(32767, 16),
 157 => to_signed(32767, 16),
 158 => to_signed(32767, 16),
 159 => to_signed(32767, 16),
 160 => to_signed(32767, 16),
 161 => to_signed(32767, 16),
 162 => to_signed(32767, 16),
 163 => to_signed(32767, 16),
 164 => to_signed(32767, 16),
 165 => to_signed(32767, 16),
 166 => to_signed(32767, 16),
 167 => to_signed(32767, 16),
 168 => to_signed(32767, 16),
 169 => to_signed(32767, 16),
 170 => to_signed(32767, 16),
 171 => to_signed(32767, 16),
 172 => to_signed(32767, 16),
 173 => to_signed(32767, 16),
 174 => to_signed(32767, 16),
 175 => to_signed(32767, 16),
 176 => to_signed(32767, 16),
 177 => to_signed(32767, 16),
 178 => to_signed(32767, 16),
 179 => to_signed(32767, 16),
 180 => to_signed(32767, 16),
 181 => to_signed(32767, 16),
 182 => to_signed(32767, 16),
 183 => to_signed(32767, 16),
 184 => to_signed(32767, 16),
 185 => to_signed(32767, 16),
 186 => to_signed(32767, 16),
 187 => to_signed(32767, 16),
 188 => to_signed(32767, 16),
 189 => to_signed(32767, 16),
 190 => to_signed(32767, 16),
 191 => to_signed(32767, 16),
 192 => to_signed(32767, 16),
 193 => to_signed(32767, 16),
 194 => to_signed(32767, 16),
 195 => to_signed(32767, 16),
 196 => to_signed(32767, 16),
 197 => to_signed(32767, 16),
 198 => to_signed(32767, 16),
 199 => to_signed(32767, 16),
 200 => to_signed(32767, 16),
 201 => to_signed(32767, 16),
 202 => to_signed(32767, 16),
 203 => to_signed(32767, 16),
 204 => to_signed(32767, 16),
 205 => to_signed(32767, 16),
 206 => to_signed(32767, 16),
 207 => to_signed(32767, 16),
 208 => to_signed(32767, 16),
 209 => to_signed(32767, 16),
 210 => to_signed(32767, 16),
 211 => to_signed(32767, 16),
 212 => to_signed(32767, 16),
 213 => to_signed(32767, 16),
 214 => to_signed(32767, 16),
 215 => to_signed(32767, 16),
 216 => to_signed(32767, 16),
 217 => to_signed(32767, 16),
 218 => to_signed(32767, 16),
 219 => to_signed(32767, 16),
 220 => to_signed(32767, 16),
 221 => to_signed(32767, 16),
 222 => to_signed(32767, 16),
 223 => to_signed(32767, 16),
 224 => to_signed(32767, 16),
 225 => to_signed(32767, 16),
 226 => to_signed(32767, 16),
 227 => to_signed(32767, 16),
 228 => to_signed(32767, 16),
 229 => to_signed(32767, 16),
 230 => to_signed(32767, 16),
 231 => to_signed(32767, 16),
 232 => to_signed(32767, 16),
 233 => to_signed(32767, 16),
 234 => to_signed(32767, 16),
 235 => to_signed(32767, 16),
 236 => to_signed(32767, 16),
 237 => to_signed(32767, 16),
 238 => to_signed(32767, 16),
 239 => to_signed(32767, 16),
 240 => to_signed(32767, 16),
 241 => to_signed(32767, 16),
 242 => to_signed(32767, 16),
 243 => to_signed(32767, 16),
 244 => to_signed(32767, 16),
 245 => to_signed(32767, 16),
 246 => to_signed(32767, 16),
 247 => to_signed(32767, 16),
 248 => to_signed(32767, 16),
 249 => to_signed(32767, 16),
 250 => to_signed(32767, 16),
 251 => to_signed(32767, 16),
 252 => to_signed(32767, 16),
 253 => to_signed(32767, 16),
 254 => to_signed(32767, 16),
 255 => to_signed(32767, 16),
 256 => to_signed(32767, 16),
 257 => to_signed(32767, 16),
 258 => to_signed(32767, 16),
 259 => to_signed(32767, 16),
 260 => to_signed(32767, 16),
 261 => to_signed(32767, 16),
 262 => to_signed(32767, 16),
 263 => to_signed(32767, 16),
 264 => to_signed(32767, 16),
 265 => to_signed(32767, 16),
 266 => to_signed(32767, 16),
 267 => to_signed(32767, 16),
 268 => to_signed(32767, 16),
 269 => to_signed(32767, 16),
 270 => to_signed(32767, 16),
 271 => to_signed(32767, 16),
 272 => to_signed(32767, 16),
 273 => to_signed(32767, 16),
 274 => to_signed(32767, 16),
 275 => to_signed(32767, 16),
 276 => to_signed(32767, 16),
 277 => to_signed(32767, 16),
 278 => to_signed(32767, 16),
 279 => to_signed(32767, 16),
 280 => to_signed(32767, 16),
 281 => to_signed(32767, 16),
 282 => to_signed(32767, 16),
 283 => to_signed(32767, 16),
 284 => to_signed(32767, 16),
 285 => to_signed(32767, 16),
 286 => to_signed(32767, 16),
 287 => to_signed(32767, 16),
 288 => to_signed(32767, 16),
 289 => to_signed(32767, 16),
 290 => to_signed(32767, 16),
 291 => to_signed(32767, 16),
 292 => to_signed(32767, 16),
 293 => to_signed(32767, 16),
 294 => to_signed(32767, 16),
 295 => to_signed(32767, 16),
 296 => to_signed(32767, 16),
 297 => to_signed(32767, 16),
 298 => to_signed(32767, 16),
 299 => to_signed(32767, 16),
 300 => to_signed(32767, 16),
 301 => to_signed(32767, 16),
 302 => to_signed(32767, 16),
 303 => to_signed(32767, 16),
 304 => to_signed(32767, 16),
 305 => to_signed(32767, 16),
 306 => to_signed(32767, 16),
 307 => to_signed(32767, 16),
 308 => to_signed(32767, 16),
 309 => to_signed(32767, 16),
 310 => to_signed(32767, 16),
 311 => to_signed(32767, 16),
 312 => to_signed(32767, 16),
 313 => to_signed(32767, 16),
 314 => to_signed(32767, 16),
 315 => to_signed(32767, 16),
 316 => to_signed(32767, 16),
 317 => to_signed(32767, 16),
 318 => to_signed(32767, 16),
 319 => to_signed(32767, 16),
 320 => to_signed(32767, 16),
 321 => to_signed(32767, 16),
 322 => to_signed(32767, 16),
 323 => to_signed(32767, 16),
 324 => to_signed(32767, 16),
 325 => to_signed(32767, 16),
 326 => to_signed(32767, 16),
 327 => to_signed(32767, 16),
 328 => to_signed(32767, 16),
 329 => to_signed(32767, 16),
 330 => to_signed(32767, 16),
 331 => to_signed(32767, 16),
 332 => to_signed(32767, 16),
 333 => to_signed(32767, 16),
 334 => to_signed(32767, 16),
 335 => to_signed(32767, 16),
 336 => to_signed(32767, 16),
 337 => to_signed(32767, 16),
 338 => to_signed(32767, 16),
 339 => to_signed(32767, 16),
 340 => to_signed(32767, 16),
 341 => to_signed(32767, 16),
 342 => to_signed(32767, 16),
 343 => to_signed(32767, 16),
 344 => to_signed(32767, 16),
 345 => to_signed(32767, 16),
 346 => to_signed(32767, 16),
 347 => to_signed(32767, 16),
 348 => to_signed(32767, 16),
 349 => to_signed(32767, 16),
 350 => to_signed(32767, 16),
 351 => to_signed(32767, 16),
 352 => to_signed(32767, 16),
 353 => to_signed(32767, 16),
 354 => to_signed(32767, 16),
 355 => to_signed(32767, 16),
 356 => to_signed(32767, 16),
 357 => to_signed(32767, 16),
 358 => to_signed(32767, 16),
 359 => to_signed(32767, 16),
 360 => to_signed(32767, 16),
 361 => to_signed(32767, 16),
 362 => to_signed(32767, 16),
 363 => to_signed(32767, 16),
 364 => to_signed(32767, 16),
 365 => to_signed(32767, 16),
 366 => to_signed(32767, 16),
 367 => to_signed(32767, 16),
 368 => to_signed(32767, 16),
 369 => to_signed(32767, 16),
 370 => to_signed(32767, 16),
 371 => to_signed(32767, 16),
 372 => to_signed(32767, 16),
 373 => to_signed(32767, 16),
 374 => to_signed(32767, 16),
 375 => to_signed(32767, 16),
 376 => to_signed(32767, 16),
 377 => to_signed(32767, 16),
 378 => to_signed(32767, 16),
 379 => to_signed(32767, 16),
 380 => to_signed(32767, 16),
 381 => to_signed(32767, 16),
 382 => to_signed(32767, 16),
 383 => to_signed(32767, 16),
 384 => to_signed(32767, 16),
 385 => to_signed(32767, 16),
 386 => to_signed(32767, 16),
 387 => to_signed(32767, 16),
 388 => to_signed(32767, 16),
 389 => to_signed(32767, 16),
 390 => to_signed(32767, 16),
 391 => to_signed(32767, 16),
 392 => to_signed(32767, 16),
 393 => to_signed(32767, 16),
 394 => to_signed(32767, 16),
 395 => to_signed(32767, 16),
 396 => to_signed(32767, 16),
 397 => to_signed(32767, 16),
 398 => to_signed(32767, 16),
 399 => to_signed(32767, 16),
 400 => to_signed(32767, 16),
 401 => to_signed(32767, 16),
 402 => to_signed(32767, 16),
 403 => to_signed(32767, 16),
 404 => to_signed(32767, 16),
 405 => to_signed(32767, 16),
 406 => to_signed(32767, 16),
 407 => to_signed(32767, 16),
 408 => to_signed(32767, 16),
 409 => to_signed(32767, 16),
 410 => to_signed(32767, 16),
 411 => to_signed(32767, 16),
 412 => to_signed(32767, 16),
 413 => to_signed(32767, 16),
 414 => to_signed(32767, 16),
 415 => to_signed(32767, 16),
 416 => to_signed(32767, 16),
 417 => to_signed(32767, 16),
 418 => to_signed(32767, 16),
 419 => to_signed(32767, 16),
 420 => to_signed(32767, 16),
 421 => to_signed(32767, 16),
 422 => to_signed(32767, 16),
 423 => to_signed(32767, 16),
 424 => to_signed(32767, 16),
 425 => to_signed(32767, 16),
 426 => to_signed(32767, 16),
 427 => to_signed(32767, 16),
 428 => to_signed(32767, 16),
 429 => to_signed(32767, 16),
 430 => to_signed(32767, 16),
 431 => to_signed(32767, 16),
 432 => to_signed(32767, 16),
 433 => to_signed(32767, 16),
 434 => to_signed(32767, 16),
 435 => to_signed(32767, 16),
 436 => to_signed(32767, 16),
 437 => to_signed(32767, 16),
 438 => to_signed(32767, 16),
 439 => to_signed(32767, 16),
 440 => to_signed(32767, 16),
 441 => to_signed(32767, 16),
 442 => to_signed(32767, 16),
 443 => to_signed(32767, 16),
 444 => to_signed(32767, 16),
 445 => to_signed(32767, 16),
 446 => to_signed(32767, 16),
 447 => to_signed(32767, 16),
 448 => to_signed(32767, 16),
 449 => to_signed(32767, 16),
 450 => to_signed(32767, 16),
 451 => to_signed(32767, 16),
 452 => to_signed(32767, 16),
 453 => to_signed(32767, 16),
 454 => to_signed(32767, 16),
 455 => to_signed(32767, 16),
 456 => to_signed(32767, 16),
 457 => to_signed(32767, 16),
 458 => to_signed(32767, 16),
 459 => to_signed(32767, 16),
 460 => to_signed(32767, 16),
 461 => to_signed(32767, 16),
 462 => to_signed(32767, 16),
 463 => to_signed(32767, 16),
 464 => to_signed(32767, 16),
 465 => to_signed(32767, 16),
 466 => to_signed(32767, 16),
 467 => to_signed(32767, 16),
 468 => to_signed(32767, 16),
 469 => to_signed(32767, 16),
 470 => to_signed(32767, 16),
 471 => to_signed(32767, 16),
 472 => to_signed(32767, 16),
 473 => to_signed(32767, 16),
 474 => to_signed(32767, 16),
 475 => to_signed(32767, 16),
 476 => to_signed(32767, 16),
 477 => to_signed(32767, 16),
 478 => to_signed(32767, 16),
 479 => to_signed(32767, 16),
 480 => to_signed(32767, 16),
 481 => to_signed(32767, 16),
 482 => to_signed(32767, 16),
 483 => to_signed(32767, 16),
 484 => to_signed(32767, 16),
 485 => to_signed(32767, 16),
 486 => to_signed(32767, 16),
 487 => to_signed(32767, 16),
 488 => to_signed(32767, 16),
 489 => to_signed(32767, 16),
 490 => to_signed(32767, 16),
 491 => to_signed(32767, 16),
 492 => to_signed(32767, 16),
 493 => to_signed(32767, 16),
 494 => to_signed(32767, 16),
 495 => to_signed(32767, 16),
 496 => to_signed(32767, 16),
 497 => to_signed(32767, 16),
 498 => to_signed(32767, 16),
 499 => to_signed(32767, 16),
 500 => to_signed(32767, 16),
 501 => to_signed(32767, 16),
 502 => to_signed(32767, 16),
 503 => to_signed(32767, 16),
 504 => to_signed(32767, 16),
 505 => to_signed(32767, 16),
 506 => to_signed(32767, 16),
 507 => to_signed(32767, 16),
 508 => to_signed(32767, 16),
 509 => to_signed(32767, 16),
 510 => to_signed(32767, 16),
 511 => to_signed(32767, 16),
 512 => to_signed(32767, 16),
 513 => to_signed(32767, 16),
 514 => to_signed(32767, 16),
 515 => to_signed(32767, 16),
 516 => to_signed(32767, 16),
 517 => to_signed(32767, 16),
 518 => to_signed(32767, 16),
 519 => to_signed(32767, 16),
 520 => to_signed(32767, 16),
 521 => to_signed(32767, 16),
 522 => to_signed(32767, 16),
 523 => to_signed(32767, 16),
 524 => to_signed(32767, 16),
 525 => to_signed(32767, 16),
 526 => to_signed(32767, 16),
 527 => to_signed(32767, 16),
 528 => to_signed(32767, 16),
 529 => to_signed(32767, 16),
 530 => to_signed(32767, 16),
 531 => to_signed(32767, 16),
 532 => to_signed(32767, 16),
 533 => to_signed(32767, 16),
 534 => to_signed(32767, 16),
 535 => to_signed(32767, 16),
 536 => to_signed(32767, 16),
 537 => to_signed(32767, 16),
 538 => to_signed(32767, 16),
 539 => to_signed(32767, 16),
 540 => to_signed(32767, 16),
 541 => to_signed(32767, 16),
 542 => to_signed(32767, 16),
 543 => to_signed(32767, 16),
 544 => to_signed(32767, 16),
 545 => to_signed(32767, 16),
 546 => to_signed(32767, 16),
 547 => to_signed(32767, 16),
 548 => to_signed(32767, 16),
 549 => to_signed(32767, 16),
 550 => to_signed(32767, 16),
 551 => to_signed(32767, 16),
 552 => to_signed(32767, 16),
 553 => to_signed(32767, 16),
 554 => to_signed(32767, 16),
 555 => to_signed(32767, 16),
 556 => to_signed(32767, 16),
 557 => to_signed(32767, 16),
 558 => to_signed(32767, 16),
 559 => to_signed(32767, 16),
 560 => to_signed(32767, 16),
 561 => to_signed(32767, 16),
 562 => to_signed(32767, 16),
 563 => to_signed(32767, 16),
 564 => to_signed(32767, 16),
 565 => to_signed(32767, 16),
 566 => to_signed(32767, 16),
 567 => to_signed(32767, 16),
 568 => to_signed(32767, 16),
 569 => to_signed(32767, 16),
 570 => to_signed(32767, 16),
 571 => to_signed(32767, 16),
 572 => to_signed(32767, 16),
 573 => to_signed(32767, 16),
 574 => to_signed(32767, 16),
 575 => to_signed(32767, 16),
 576 => to_signed(32767, 16),
 577 => to_signed(32767, 16),
 578 => to_signed(32767, 16),
 579 => to_signed(32767, 16),
 580 => to_signed(32767, 16),
 581 => to_signed(32767, 16),
 582 => to_signed(32767, 16),
 583 => to_signed(32767, 16),
 584 => to_signed(32767, 16),
 585 => to_signed(32767, 16),
 586 => to_signed(32767, 16),
 587 => to_signed(32767, 16),
 588 => to_signed(32767, 16),
 589 => to_signed(32767, 16),
 590 => to_signed(32767, 16),
 591 => to_signed(32767, 16),
 592 => to_signed(32767, 16),
 593 => to_signed(32767, 16),
 594 => to_signed(32767, 16),
 595 => to_signed(32767, 16),
 596 => to_signed(32767, 16),
 597 => to_signed(32767, 16),
 598 => to_signed(32767, 16),
 599 => to_signed(32767, 16),
 600 => to_signed(32767, 16),
 601 => to_signed(32767, 16),
 602 => to_signed(32767, 16),
 603 => to_signed(32767, 16),
 604 => to_signed(32767, 16),
 605 => to_signed(32767, 16),
 606 => to_signed(32767, 16),
 607 => to_signed(32767, 16),
 608 => to_signed(32767, 16),
 609 => to_signed(32767, 16),
 610 => to_signed(32767, 16),
 611 => to_signed(32767, 16),
 612 => to_signed(32767, 16),
 613 => to_signed(32767, 16),
 614 => to_signed(32767, 16),
 615 => to_signed(32767, 16),
 616 => to_signed(32767, 16),
 617 => to_signed(32767, 16),
 618 => to_signed(32767, 16),
 619 => to_signed(32767, 16),
 620 => to_signed(32767, 16),
 621 => to_signed(32767, 16),
 622 => to_signed(32767, 16),
 623 => to_signed(32767, 16),
 624 => to_signed(32767, 16),
 625 => to_signed(32767, 16),
 626 => to_signed(32767, 16),
 627 => to_signed(32767, 16),
 628 => to_signed(32767, 16),
 629 => to_signed(32767, 16),
 630 => to_signed(32767, 16),
 631 => to_signed(32767, 16),
 632 => to_signed(32767, 16),
 633 => to_signed(32767, 16),
 634 => to_signed(32767, 16),
 635 => to_signed(32767, 16),
 636 => to_signed(32767, 16),
 637 => to_signed(32767, 16),
 638 => to_signed(32767, 16),
 639 => to_signed(32767, 16),
 640 => to_signed(32767, 16),
 641 => to_signed(32767, 16),
 642 => to_signed(32767, 16),
 643 => to_signed(32767, 16),
 644 => to_signed(32767, 16),
 645 => to_signed(32767, 16),
 646 => to_signed(32767, 16),
 647 => to_signed(32767, 16),
 648 => to_signed(32767, 16),
 649 => to_signed(32767, 16),
 650 => to_signed(32767, 16),
 651 => to_signed(32767, 16),
 652 => to_signed(32767, 16),
 653 => to_signed(32767, 16),
 654 => to_signed(32767, 16),
 655 => to_signed(32767, 16),
 656 => to_signed(32767, 16),
 657 => to_signed(32767, 16),
 658 => to_signed(32767, 16),
 659 => to_signed(32767, 16),
 660 => to_signed(32767, 16),
 661 => to_signed(32767, 16),
 662 => to_signed(32767, 16),
 663 => to_signed(32767, 16),
 664 => to_signed(32767, 16),
 665 => to_signed(32767, 16),
 666 => to_signed(32767, 16),
 667 => to_signed(32767, 16),
 668 => to_signed(32767, 16),
 669 => to_signed(32767, 16),
 670 => to_signed(32767, 16),
 671 => to_signed(32767, 16),
 672 => to_signed(32767, 16),
 673 => to_signed(32767, 16),
 674 => to_signed(32767, 16),
 675 => to_signed(32767, 16),
 676 => to_signed(32767, 16),
 677 => to_signed(32767, 16),
 678 => to_signed(32767, 16),
 679 => to_signed(32767, 16),
 680 => to_signed(32767, 16),
 681 => to_signed(32767, 16),
 682 => to_signed(32767, 16),
 683 => to_signed(32767, 16),
 684 => to_signed(32767, 16),
 685 => to_signed(32767, 16),
 686 => to_signed(32767, 16),
 687 => to_signed(32767, 16),
 688 => to_signed(32767, 16),
 689 => to_signed(32767, 16),
 690 => to_signed(32767, 16),
 691 => to_signed(32767, 16),
 692 => to_signed(32767, 16),
 693 => to_signed(32767, 16),
 694 => to_signed(32767, 16),
 695 => to_signed(32767, 16),
 696 => to_signed(32767, 16),
 697 => to_signed(32767, 16),
 698 => to_signed(32767, 16),
 699 => to_signed(32767, 16),
 700 => to_signed(32767, 16),
 701 => to_signed(32767, 16),
 702 => to_signed(32767, 16),
 703 => to_signed(32767, 16),
 704 => to_signed(32767, 16),
 705 => to_signed(32767, 16),
 706 => to_signed(32767, 16),
 707 => to_signed(32767, 16),
 708 => to_signed(32767, 16),
 709 => to_signed(32767, 16),
 710 => to_signed(32767, 16),
 711 => to_signed(32767, 16),
 712 => to_signed(32767, 16),
 713 => to_signed(32767, 16),
 714 => to_signed(32767, 16),
 715 => to_signed(32767, 16),
 716 => to_signed(32767, 16),
 717 => to_signed(32767, 16),
 718 => to_signed(32767, 16),
 719 => to_signed(32767, 16),
 720 => to_signed(32767, 16),
 721 => to_signed(32767, 16),
 722 => to_signed(32767, 16),
 723 => to_signed(32767, 16),
 724 => to_signed(32767, 16),
 725 => to_signed(32767, 16),
 726 => to_signed(32767, 16),
 727 => to_signed(32767, 16),
 728 => to_signed(32767, 16),
 729 => to_signed(32767, 16),
 730 => to_signed(32767, 16),
 731 => to_signed(32767, 16),
 732 => to_signed(32767, 16),
 733 => to_signed(32767, 16),
 734 => to_signed(32767, 16),
 735 => to_signed(32767, 16),
 736 => to_signed(32767, 16),
 737 => to_signed(32767, 16),
 738 => to_signed(32767, 16),
 739 => to_signed(32767, 16),
 740 => to_signed(32767, 16),
 741 => to_signed(32767, 16),
 742 => to_signed(32767, 16),
 743 => to_signed(32767, 16),
 744 => to_signed(32767, 16),
 745 => to_signed(32767, 16),
 746 => to_signed(32767, 16),
 747 => to_signed(32767, 16),
 748 => to_signed(32767, 16),
 749 => to_signed(32767, 16),
 750 => to_signed(32767, 16),
 751 => to_signed(32767, 16),
 752 => to_signed(32767, 16),
 753 => to_signed(32767, 16),
 754 => to_signed(32767, 16),
 755 => to_signed(32767, 16),
 756 => to_signed(32767, 16),
 757 => to_signed(32767, 16),
 758 => to_signed(32767, 16),
 759 => to_signed(32767, 16),
 760 => to_signed(32767, 16),
 761 => to_signed(32767, 16),
 762 => to_signed(32767, 16),
 763 => to_signed(32767, 16),
 764 => to_signed(32767, 16),
 765 => to_signed(32767, 16),
 766 => to_signed(32767, 16),
 767 => to_signed(32767, 16),
 768 => to_signed(32767, 16),
 769 => to_signed(32767, 16),
 770 => to_signed(32767, 16),
 771 => to_signed(32767, 16),
 772 => to_signed(32767, 16),
 773 => to_signed(32767, 16),
 774 => to_signed(32767, 16),
 775 => to_signed(32767, 16),
 776 => to_signed(32767, 16),
 777 => to_signed(32767, 16),
 778 => to_signed(32767, 16),
 779 => to_signed(32767, 16),
 780 => to_signed(32767, 16),
 781 => to_signed(32767, 16),
 782 => to_signed(32767, 16),
 783 => to_signed(32767, 16),
 784 => to_signed(32767, 16),
 785 => to_signed(32767, 16),
 786 => to_signed(32767, 16),
 787 => to_signed(32767, 16),
 788 => to_signed(32767, 16),
 789 => to_signed(32767, 16),
 790 => to_signed(32767, 16),
 791 => to_signed(32767, 16),
 792 => to_signed(32767, 16),
 793 => to_signed(32767, 16),
 794 => to_signed(32767, 16),
 795 => to_signed(32767, 16),
 796 => to_signed(32767, 16),
 797 => to_signed(32767, 16),
 798 => to_signed(32767, 16),
 799 => to_signed(32767, 16),
 800 => to_signed(32767, 16),
 801 => to_signed(32767, 16),
 802 => to_signed(32767, 16),
 803 => to_signed(32767, 16),
 804 => to_signed(32767, 16),
 805 => to_signed(32767, 16),
 806 => to_signed(32767, 16),
 807 => to_signed(32767, 16),
 808 => to_signed(32767, 16),
 809 => to_signed(32767, 16),
 810 => to_signed(32767, 16),
 811 => to_signed(32767, 16),
 812 => to_signed(32767, 16),
 813 => to_signed(32767, 16),
 814 => to_signed(32767, 16),
 815 => to_signed(32767, 16),
 816 => to_signed(32767, 16),
 817 => to_signed(32767, 16),
 818 => to_signed(32767, 16),
 819 => to_signed(32767, 16),
 820 => to_signed(32767, 16),
 821 => to_signed(32767, 16),
 822 => to_signed(32767, 16),
 823 => to_signed(32767, 16),
 824 => to_signed(32767, 16),
 825 => to_signed(32767, 16),
 826 => to_signed(32767, 16),
 827 => to_signed(32767, 16),
 828 => to_signed(32767, 16),
 829 => to_signed(32767, 16),
 830 => to_signed(32767, 16),
 831 => to_signed(32767, 16),
 832 => to_signed(32767, 16),
 833 => to_signed(32767, 16),
 834 => to_signed(32767, 16),
 835 => to_signed(32767, 16),
 836 => to_signed(32767, 16),
 837 => to_signed(32767, 16),
 838 => to_signed(32767, 16),
 839 => to_signed(32767, 16),
 840 => to_signed(32767, 16),
 841 => to_signed(32767, 16),
 842 => to_signed(32767, 16),
 843 => to_signed(32767, 16),
 844 => to_signed(32767, 16),
 845 => to_signed(32767, 16),
 846 => to_signed(32767, 16),
 847 => to_signed(32767, 16),
 848 => to_signed(32767, 16),
 849 => to_signed(32767, 16),
 850 => to_signed(32767, 16),
 851 => to_signed(32767, 16),
 852 => to_signed(32767, 16),
 853 => to_signed(32767, 16),
 854 => to_signed(32767, 16),
 855 => to_signed(32767, 16),
 856 => to_signed(32767, 16),
 857 => to_signed(32767, 16),
 858 => to_signed(32767, 16),
 859 => to_signed(32767, 16),
 860 => to_signed(32767, 16),
 861 => to_signed(32767, 16),
 862 => to_signed(32767, 16),
 863 => to_signed(32767, 16),
 864 => to_signed(32767, 16),
 865 => to_signed(32767, 16),
 866 => to_signed(32767, 16),
 867 => to_signed(32767, 16),
 868 => to_signed(32767, 16),
 869 => to_signed(32767, 16),
 870 => to_signed(32767, 16),
 871 => to_signed(32767, 16),
 872 => to_signed(32767, 16),
 873 => to_signed(32767, 16),
 874 => to_signed(32767, 16),
 875 => to_signed(32767, 16),
 876 => to_signed(32767, 16),
 877 => to_signed(32767, 16),
 878 => to_signed(32767, 16),
 879 => to_signed(32767, 16),
 880 => to_signed(32767, 16),
 881 => to_signed(32767, 16),
 882 => to_signed(32767, 16),
 883 => to_signed(32767, 16),
 884 => to_signed(32767, 16),
 885 => to_signed(32767, 16),
 886 => to_signed(32767, 16),
 887 => to_signed(32767, 16),
 888 => to_signed(32767, 16),
 889 => to_signed(32767, 16),
 890 => to_signed(32767, 16),
 891 => to_signed(32767, 16),
 892 => to_signed(32767, 16),
 893 => to_signed(32767, 16),
 894 => to_signed(32767, 16),
 895 => to_signed(32767, 16),
 896 => to_signed(32767, 16),
 897 => to_signed(32767, 16),
 898 => to_signed(32767, 16),
 899 => to_signed(32767, 16));

type DATA_OUT_ARRAY_T is array (natural range <>) of signed(17 downto 0);
constant DATA_OUT_ARRAY : DATA_OUT_ARRAY_T(0 to 899) :=
(0 => to_signed(32047, 18),
 1 => to_signed(30624, 18),
 2 => to_signed(29232, 18),
 3 => to_signed(27873, 18),
 4 => to_signed(26547, 18),
 5 => to_signed(25253, 18),
 6 => to_signed(23990, 18),
 7 => to_signed(22760, 18),
 8 => to_signed(21561, 18),
 9 => to_signed(20394, 18),
 10 => to_signed(19257, 18),
 11 => to_signed(18152, 18),
 12 => to_signed(17077, 18),
 13 => to_signed(16033, 18),
 14 => to_signed(15018, 18),
 15 => to_signed(14034, 18),
 16 => to_signed(13078, 18),
 17 => to_signed(12152, 18),
 18 => to_signed(11254, 18),
 19 => to_signed(10385, 18),
 20 => to_signed(9543, 18),
 21 => to_signed(8729, 18),
 22 => to_signed(7941, 18),
 23 => to_signed(7181, 18),
 24 => to_signed(6446, 18),
 25 => to_signed(5738, 18),
 26 => to_signed(5054, 18),
 27 => to_signed(4396, 18),
 28 => to_signed(3761, 18),
 29 => to_signed(3151, 18),
 30 => to_signed(2564, 18),
 31 => to_signed(2001, 18),
 32 => to_signed(1459, 18),
 33 => to_signed(941, 18),
 34 => to_signed(442, 18),
 35 => to_signed(-33, 18),
 36 => to_signed(-489, 18),
 37 => to_signed(-924, 18),
 38 => to_signed(-1340, 18),
 39 => to_signed(-1735, 18),
 40 => to_signed(-2113, 18),
 41 => to_signed(-2471, 18),
 42 => to_signed(-2812, 18),
 43 => to_signed(-3135, 18),
 44 => to_signed(-3442, 18),
 45 => to_signed(-3731, 18),
 46 => to_signed(-4005, 18),
 47 => to_signed(-4262, 18),
 48 => to_signed(-4505, 18),
 49 => to_signed(-4732, 18),
 50 => to_signed(-4946, 18),
 51 => to_signed(-5144, 18),
 52 => to_signed(-5330, 18),
 53 => to_signed(-5502, 18),
 54 => to_signed(-5662, 18),
 55 => to_signed(-5809, 18),
 56 => to_signed(-5944, 18),
 57 => to_signed(-6068, 18),
 58 => to_signed(-6181, 18),
 59 => to_signed(-6282, 18),
 60 => to_signed(-6373, 18),
 61 => to_signed(-6454, 18),
 62 => to_signed(-6526, 18),
 63 => to_signed(-6588, 18),
 64 => to_signed(-6641, 18),
 65 => to_signed(-6685, 18),
 66 => to_signed(-6721, 18),
 67 => to_signed(-6749, 18),
 68 => to_signed(-6769, 18),
 69 => to_signed(-6782, 18),
 70 => to_signed(-6788, 18),
 71 => to_signed(-6787, 18),
 72 => to_signed(-6780, 18),
 73 => to_signed(-6766, 18),
 74 => to_signed(-6747, 18),
 75 => to_signed(-6722, 18),
 76 => to_signed(-6691, 18),
 77 => to_signed(-6656, 18),
 78 => to_signed(-6615, 18),
 79 => to_signed(-6570, 18),
 80 => to_signed(-6521, 18),
 81 => to_signed(-6467, 18),
 82 => to_signed(-6410, 18),
 83 => to_signed(-6349, 18),
 84 => to_signed(-6285, 18),
 85 => to_signed(-6217, 18),
 86 => to_signed(-6147, 18),
 87 => to_signed(-6073, 18),
 88 => to_signed(-5997, 18),
 89 => to_signed(-5918, 18),
 90 => to_signed(-5838, 18),
 91 => to_signed(-5754, 18),
 92 => to_signed(-5670, 18),
 93 => to_signed(-5583, 18),
 94 => to_signed(-5495, 18),
 95 => to_signed(-5405, 18),
 96 => to_signed(-5314, 18),
 97 => to_signed(-5222, 18),
 98 => to_signed(-5129, 18),
 99 => to_signed(-5035, 18),
 100 => to_signed(-4941, 18),
 101 => to_signed(-4845, 18),
 102 => to_signed(-4749, 18),
 103 => to_signed(-4653, 18),
 104 => to_signed(-4557, 18),
 105 => to_signed(-4459, 18),
 106 => to_signed(-4363, 18),
 107 => to_signed(-4266, 18),
 108 => to_signed(-4170, 18),
 109 => to_signed(-4073, 18),
 110 => to_signed(-3977, 18),
 111 => to_signed(-3881, 18),
 112 => to_signed(-3786, 18),
 113 => to_signed(-3691, 18),
 114 => to_signed(-3597, 18),
 115 => to_signed(-3503, 18),
 116 => to_signed(-3410, 18),
 117 => to_signed(-3318, 18),
 118 => to_signed(-3227, 18),
 119 => to_signed(-3136, 18),
 120 => to_signed(-3047, 18),
 121 => to_signed(-2958, 18),
 122 => to_signed(-2871, 18),
 123 => to_signed(-2784, 18),
 124 => to_signed(-2699, 18),
 125 => to_signed(-2615, 18),
 126 => to_signed(-2531, 18),
 127 => to_signed(-2450, 18),
 128 => to_signed(-2368, 18),
 129 => to_signed(-2289, 18),
 130 => to_signed(-2211, 18),
 131 => to_signed(-2134, 18),
 132 => to_signed(-2058, 18),
 133 => to_signed(-1984, 18),
 134 => to_signed(-1911, 18),
 135 => to_signed(-1840, 18),
 136 => to_signed(-1769, 18),
 137 => to_signed(-1700, 18),
 138 => to_signed(-1632, 18),
 139 => to_signed(-1566, 18),
 140 => to_signed(-1501, 18),
 141 => to_signed(-1438, 18),
 142 => to_signed(-1375, 18),
 143 => to_signed(-1315, 18),
 144 => to_signed(-1255, 18),
 145 => to_signed(-1198, 18),
 146 => to_signed(-1141, 18),
 147 => to_signed(-1086, 18),
 148 => to_signed(-1032, 18),
 149 => to_signed(-980, 18),
 150 => to_signed(-928, 18),
 151 => to_signed(-879, 18),
 152 => to_signed(-830, 18),
 153 => to_signed(-783, 18),
 154 => to_signed(-736, 18),
 155 => to_signed(-692, 18),
 156 => to_signed(-648, 18),
 157 => to_signed(-607, 18),
 158 => to_signed(-565, 18),
 159 => to_signed(-527, 18),
 160 => to_signed(-487, 18),
 161 => to_signed(-451, 18),
 162 => to_signed(-414, 18),
 163 => to_signed(-380, 18),
 164 => to_signed(-346, 18),
 165 => to_signed(-314, 18),
 166 => to_signed(-282, 18),
 167 => to_signed(-252, 18),
 168 => to_signed(-222, 18),
 169 => to_signed(-195, 18),
 170 => to_signed(-166, 18),
 171 => to_signed(-142, 18),
 172 => to_signed(-115, 18),
 173 => to_signed(-93, 18),
 174 => to_signed(-68, 18),
 175 => to_signed(-47, 18),
 176 => to_signed(-24, 18),
 177 => to_signed(-5, 18),
 178 => to_signed(16, 18),
 179 => to_signed(33, 18),
 180 => to_signed(53, 18),
 181 => to_signed(68, 18),
 182 => to_signed(86, 18),
 183 => to_signed(99, 18),
 184 => to_signed(116, 18),
 185 => to_signed(128, 18),
 186 => to_signed(143, 18),
 187 => to_signed(153, 18),
 188 => to_signed(167, 18),
 189 => to_signed(176, 18),
 190 => to_signed(189, 18),
 191 => to_signed(197, 18),
 192 => to_signed(208, 18),
 193 => to_signed(214, 18),
 194 => to_signed(225, 18),
 195 => to_signed(230, 18),
 196 => to_signed(239, 18),
 197 => to_signed(243, 18),
 198 => to_signed(251, 18),
 199 => to_signed(255, 18),
 200 => to_signed(261, 18),
 201 => to_signed(264, 18),
 202 => to_signed(270, 18),
 203 => to_signed(272, 18),
 204 => to_signed(276, 18),
 205 => to_signed(278, 18),
 206 => to_signed(281, 18),
 207 => to_signed(282, 18),
 208 => to_signed(285, 18),
 209 => to_signed(285, 18),
 210 => to_signed(287, 18),
 211 => to_signed(286, 18),
 212 => to_signed(288, 18),
 213 => to_signed(287, 18),
 214 => to_signed(288, 18),
 215 => to_signed(286, 18),
 216 => to_signed(287, 18),
 217 => to_signed(284, 18),
 218 => to_signed(285, 18),
 219 => to_signed(282, 18),
 220 => to_signed(282, 18),
 221 => to_signed(278, 18),
 222 => to_signed(278, 18),
 223 => to_signed(274, 18),
 224 => to_signed(273, 18),
 225 => to_signed(269, 18),
 226 => to_signed(268, 18),
 227 => to_signed(264, 18),
 228 => to_signed(262, 18),
 229 => to_signed(258, 18),
 230 => to_signed(256, 18),
 231 => to_signed(251, 18),
 232 => to_signed(249, 18),
 233 => to_signed(244, 18),
 234 => to_signed(242, 18),
 235 => to_signed(237, 18),
 236 => to_signed(234, 18),
 237 => to_signed(230, 18),
 238 => to_signed(227, 18),
 239 => to_signed(222, 18),
 240 => to_signed(219, 18),
 241 => to_signed(214, 18),
 242 => to_signed(211, 18),
 243 => to_signed(206, 18),
 244 => to_signed(202, 18),
 245 => to_signed(198, 18),
 246 => to_signed(194, 18),
 247 => to_signed(190, 18),
 248 => to_signed(186, 18),
 249 => to_signed(182, 18),
 250 => to_signed(178, 18),
 251 => to_signed(174, 18),
 252 => to_signed(169, 18),
 253 => to_signed(166, 18),
 254 => to_signed(161, 18),
 255 => to_signed(158, 18),
 256 => to_signed(153, 18),
 257 => to_signed(150, 18),
 258 => to_signed(145, 18),
 259 => to_signed(143, 18),
 260 => to_signed(137, 18),
 261 => to_signed(135, 18),
 262 => to_signed(129, 18),
 263 => to_signed(127, 18),
 264 => to_signed(122, 18),
 265 => to_signed(120, 18),
 266 => to_signed(115, 18),
 267 => to_signed(113, 18),
 268 => to_signed(107, 18),
 269 => to_signed(106, 18),
 270 => to_signed(101, 18),
 271 => to_signed(99, 18),
 272 => to_signed(94, 18),
 273 => to_signed(92, 18),
 274 => to_signed(87, 18),
 275 => to_signed(86, 18),
 276 => to_signed(81, 18),
 277 => to_signed(80, 18),
 278 => to_signed(75, 18),
 279 => to_signed(74, 18),
 280 => to_signed(69, 18),
 281 => to_signed(68, 18),
 282 => to_signed(63, 18),
 283 => to_signed(63, 18),
 284 => to_signed(58, 18),
 285 => to_signed(58, 18),
 286 => to_signed(53, 18),
 287 => to_signed(53, 18),
 288 => to_signed(48, 18),
 289 => to_signed(48, 18),
 290 => to_signed(43, 18),
 291 => to_signed(43, 18),
 292 => to_signed(39, 18),
 293 => to_signed(39, 18),
 294 => to_signed(35, 18),
 295 => to_signed(35, 18),
 296 => to_signed(31, 18),
 297 => to_signed(31, 18),
 298 => to_signed(27, 18),
 299 => to_signed(27, 18),
 300 => to_signed(24, 18),
 301 => to_signed(24, 18),
 302 => to_signed(21, 18),
 303 => to_signed(20, 18),
 304 => to_signed(18, 18),
 305 => to_signed(17, 18),
 306 => to_signed(15, 18),
 307 => to_signed(14, 18),
 308 => to_signed(12, 18),
 309 => to_signed(11, 18),
 310 => to_signed(10, 18),
 311 => to_signed(9, 18),
 312 => to_signed(8, 18),
 313 => to_signed(6, 18),
 314 => to_signed(5, 18),
 315 => to_signed(4, 18),
 316 => to_signed(4, 18),
 317 => to_signed(2, 18),
 318 => to_signed(2, 18),
 319 => to_signed(0, 18),
 320 => to_signed(0, 18),
 321 => to_signed(-2, 18),
 322 => to_signed(-1, 18),
 323 => to_signed(-3, 18),
 324 => to_signed(-3, 18),
 325 => to_signed(-5, 18),
 326 => to_signed(-4, 18),
 327 => to_signed(-6, 18),
 328 => to_signed(-5, 18),
 329 => to_signed(-7, 18),
 330 => to_signed(-6, 18),
 331 => to_signed(-8, 18),
 332 => to_signed(-7, 18),
 333 => to_signed(-9, 18),
 334 => to_signed(-8, 18),
 335 => to_signed(-10, 18),
 336 => to_signed(-8, 18),
 337 => to_signed(-11, 18),
 338 => to_signed(-9, 18),
 339 => to_signed(-11, 18),
 340 => to_signed(-10, 18),
 341 => to_signed(-11, 18),
 342 => to_signed(-10, 18),
 343 => to_signed(-12, 18),
 344 => to_signed(-11, 18),
 345 => to_signed(-12, 18),
 346 => to_signed(-11, 18),
 347 => to_signed(-12, 18),
 348 => to_signed(-11, 18),
 349 => to_signed(-12, 18),
 350 => to_signed(-12, 18),
 351 => to_signed(-12, 18),
 352 => to_signed(-12, 18),
 353 => to_signed(-12, 18),
 354 => to_signed(-12, 18),
 355 => to_signed(-12, 18),
 356 => to_signed(-12, 18),
 357 => to_signed(-12, 18),
 358 => to_signed(-12, 18),
 359 => to_signed(-12, 18),
 360 => to_signed(-12, 18),
 361 => to_signed(-12, 18),
 362 => to_signed(-12, 18),
 363 => to_signed(-12, 18),
 364 => to_signed(-12, 18),
 365 => to_signed(-12, 18),
 366 => to_signed(-12, 18),
 367 => to_signed(-11, 18),
 368 => to_signed(-11, 18),
 369 => to_signed(-11, 18),
 370 => to_signed(-11, 18),
 371 => to_signed(-11, 18),
 372 => to_signed(-11, 18),
 373 => to_signed(-11, 18),
 374 => to_signed(-10, 18),
 375 => to_signed(-10, 18),
 376 => to_signed(-10, 18),
 377 => to_signed(-10, 18),
 378 => to_signed(-10, 18),
 379 => to_signed(-10, 18),
 380 => to_signed(-10, 18),
 381 => to_signed(-10, 18),
 382 => to_signed(-9, 18),
 383 => to_signed(-9, 18),
 384 => to_signed(-9, 18),
 385 => to_signed(-9, 18),
 386 => to_signed(-9, 18),
 387 => to_signed(-8, 18),
 388 => to_signed(-8, 18),
 389 => to_signed(-8, 18),
 390 => to_signed(-8, 18),
 391 => to_signed(-8, 18),
 392 => to_signed(-8, 18),
 393 => to_signed(-7, 18),
 394 => to_signed(-7, 18),
 395 => to_signed(-7, 18),
 396 => to_signed(-7, 18),
 397 => to_signed(-7, 18),
 398 => to_signed(-7, 18),
 399 => to_signed(-6, 18),
 400 => to_signed(-6, 18),
 401 => to_signed(-6, 18),
 402 => to_signed(-6, 18),
 403 => to_signed(-5, 18),
 404 => to_signed(-6, 18),
 405 => to_signed(-5, 18),
 406 => to_signed(-5, 18),
 407 => to_signed(-5, 18),
 408 => to_signed(-5, 18),
 409 => to_signed(-5, 18),
 410 => to_signed(-5, 18),
 411 => to_signed(-4, 18),
 412 => to_signed(-5, 18),
 413 => to_signed(-4, 18),
 414 => to_signed(-4, 18),
 415 => to_signed(-4, 18),
 416 => to_signed(-4, 18),
 417 => to_signed(-3, 18),
 418 => to_signed(-4, 18),
 419 => to_signed(-3, 18),
 420 => to_signed(-3, 18),
 421 => to_signed(-3, 18),
 422 => to_signed(-3, 18),
 423 => to_signed(-3, 18),
 424 => to_signed(-3, 18),
 425 => to_signed(-3, 18),
 426 => to_signed(-2, 18),
 427 => to_signed(-3, 18),
 428 => to_signed(-2, 18),
 429 => to_signed(-2, 18),
 430 => to_signed(-2, 18),
 431 => to_signed(-2, 18),
 432 => to_signed(-2, 18),
 433 => to_signed(-2, 18),
 434 => to_signed(-2, 18),
 435 => to_signed(-2, 18),
 436 => to_signed(-1, 18),
 437 => to_signed(-2, 18),
 438 => to_signed(-1, 18),
 439 => to_signed(-1, 18),
 440 => to_signed(-1, 18),
 441 => to_signed(-1, 18),
 442 => to_signed(-1, 18),
 443 => to_signed(-1, 18),
 444 => to_signed(-1, 18),
 445 => to_signed(-1, 18),
 446 => to_signed(0, 18),
 447 => to_signed(-1, 18),
 448 => to_signed(0, 18),
 449 => to_signed(-1, 18),
 450 => to_signed(0, 18),
 451 => to_signed(-1, 18),
 452 => to_signed(0, 18),
 453 => to_signed(-1, 18),
 454 => to_signed(0, 18),
 455 => to_signed(-1, 18),
 456 => to_signed(0, 18),
 457 => to_signed(-1, 18),
 458 => to_signed(0, 18),
 459 => to_signed(0, 18),
 460 => to_signed(0, 18),
 461 => to_signed(0, 18),
 462 => to_signed(0, 18),
 463 => to_signed(0, 18),
 464 => to_signed(1, 18),
 465 => to_signed(0, 18),
 466 => to_signed(1, 18),
 467 => to_signed(0, 18),
 468 => to_signed(1, 18),
 469 => to_signed(0, 18),
 470 => to_signed(1, 18),
 471 => to_signed(0, 18),
 472 => to_signed(1, 18),
 473 => to_signed(0, 18),
 474 => to_signed(1, 18),
 475 => to_signed(0, 18),
 476 => to_signed(1, 18),
 477 => to_signed(0, 18),
 478 => to_signed(1, 18),
 479 => to_signed(0, 18),
 480 => to_signed(1, 18),
 481 => to_signed(0, 18),
 482 => to_signed(1, 18),
 483 => to_signed(0, 18),
 484 => to_signed(1, 18),
 485 => to_signed(0, 18),
 486 => to_signed(1, 18),
 487 => to_signed(0, 18),
 488 => to_signed(1, 18),
 489 => to_signed(0, 18),
 490 => to_signed(1, 18),
 491 => to_signed(1, 18),
 492 => to_signed(0, 18),
 493 => to_signed(1, 18),
 494 => to_signed(0, 18),
 495 => to_signed(1, 18),
 496 => to_signed(0, 18),
 497 => to_signed(1, 18),
 498 => to_signed(0, 18),
 499 => to_signed(1, 18),
 500 => to_signed(0, 18),
 501 => to_signed(1, 18),
 502 => to_signed(0, 18),
 503 => to_signed(1, 18),
 504 => to_signed(0, 18),
 505 => to_signed(1, 18),
 506 => to_signed(0, 18),
 507 => to_signed(1, 18),
 508 => to_signed(0, 18),
 509 => to_signed(1, 18),
 510 => to_signed(0, 18),
 511 => to_signed(1, 18),
 512 => to_signed(0, 18),
 513 => to_signed(1, 18),
 514 => to_signed(0, 18),
 515 => to_signed(1, 18),
 516 => to_signed(0, 18),
 517 => to_signed(1, 18),
 518 => to_signed(0, 18),
 519 => to_signed(1, 18),
 520 => to_signed(0, 18),
 521 => to_signed(1, 18),
 522 => to_signed(0, 18),
 523 => to_signed(1, 18),
 524 => to_signed(0, 18),
 525 => to_signed(1, 18),
 526 => to_signed(0, 18),
 527 => to_signed(1, 18),
 528 => to_signed(0, 18),
 529 => to_signed(1, 18),
 530 => to_signed(0, 18),
 531 => to_signed(1, 18),
 532 => to_signed(0, 18),
 533 => to_signed(1, 18),
 534 => to_signed(0, 18),
 535 => to_signed(1, 18),
 536 => to_signed(0, 18),
 537 => to_signed(1, 18),
 538 => to_signed(0, 18),
 539 => to_signed(1, 18),
 540 => to_signed(0, 18),
 541 => to_signed(1, 18),
 542 => to_signed(0, 18),
 543 => to_signed(1, 18),
 544 => to_signed(0, 18),
 545 => to_signed(1, 18),
 546 => to_signed(0, 18),
 547 => to_signed(1, 18),
 548 => to_signed(0, 18),
 549 => to_signed(1, 18),
 550 => to_signed(0, 18),
 551 => to_signed(1, 18),
 552 => to_signed(0, 18),
 553 => to_signed(1, 18),
 554 => to_signed(0, 18),
 555 => to_signed(1, 18),
 556 => to_signed(0, 18),
 557 => to_signed(1, 18),
 558 => to_signed(0, 18),
 559 => to_signed(1, 18),
 560 => to_signed(0, 18),
 561 => to_signed(1, 18),
 562 => to_signed(0, 18),
 563 => to_signed(0, 18),
 564 => to_signed(0, 18),
 565 => to_signed(0, 18),
 566 => to_signed(0, 18),
 567 => to_signed(0, 18),
 568 => to_signed(0, 18),
 569 => to_signed(0, 18),
 570 => to_signed(0, 18),
 571 => to_signed(0, 18),
 572 => to_signed(0, 18),
 573 => to_signed(0, 18),
 574 => to_signed(0, 18),
 575 => to_signed(0, 18),
 576 => to_signed(0, 18),
 577 => to_signed(0, 18),
 578 => to_signed(0, 18),
 579 => to_signed(0, 18),
 580 => to_signed(0, 18),
 581 => to_signed(0, 18),
 582 => to_signed(0, 18),
 583 => to_signed(0, 18),
 584 => to_signed(0, 18),
 585 => to_signed(0, 18),
 586 => to_signed(0, 18),
 587 => to_signed(0, 18),
 588 => to_signed(0, 18),
 589 => to_signed(0, 18),
 590 => to_signed(0, 18),
 591 => to_signed(0, 18),
 592 => to_signed(0, 18),
 593 => to_signed(0, 18),
 594 => to_signed(0, 18),
 595 => to_signed(0, 18),
 596 => to_signed(0, 18),
 597 => to_signed(0, 18),
 598 => to_signed(0, 18),
 599 => to_signed(0, 18),
 600 => to_signed(0, 18),
 601 => to_signed(0, 18),
 602 => to_signed(0, 18),
 603 => to_signed(0, 18),
 604 => to_signed(0, 18),
 605 => to_signed(0, 18),
 606 => to_signed(0, 18),
 607 => to_signed(0, 18),
 608 => to_signed(0, 18),
 609 => to_signed(0, 18),
 610 => to_signed(0, 18),
 611 => to_signed(0, 18),
 612 => to_signed(0, 18),
 613 => to_signed(0, 18),
 614 => to_signed(0, 18),
 615 => to_signed(0, 18),
 616 => to_signed(0, 18),
 617 => to_signed(0, 18),
 618 => to_signed(0, 18),
 619 => to_signed(0, 18),
 620 => to_signed(0, 18),
 621 => to_signed(0, 18),
 622 => to_signed(0, 18),
 623 => to_signed(0, 18),
 624 => to_signed(0, 18),
 625 => to_signed(0, 18),
 626 => to_signed(0, 18),
 627 => to_signed(0, 18),
 628 => to_signed(0, 18),
 629 => to_signed(0, 18),
 630 => to_signed(0, 18),
 631 => to_signed(0, 18),
 632 => to_signed(0, 18),
 633 => to_signed(0, 18),
 634 => to_signed(0, 18),
 635 => to_signed(0, 18),
 636 => to_signed(0, 18),
 637 => to_signed(0, 18),
 638 => to_signed(0, 18),
 639 => to_signed(0, 18),
 640 => to_signed(0, 18),
 641 => to_signed(0, 18),
 642 => to_signed(0, 18),
 643 => to_signed(0, 18),
 644 => to_signed(0, 18),
 645 => to_signed(0, 18),
 646 => to_signed(0, 18),
 647 => to_signed(0, 18),
 648 => to_signed(0, 18),
 649 => to_signed(0, 18),
 650 => to_signed(0, 18),
 651 => to_signed(0, 18),
 652 => to_signed(0, 18),
 653 => to_signed(0, 18),
 654 => to_signed(0, 18),
 655 => to_signed(0, 18),
 656 => to_signed(0, 18),
 657 => to_signed(0, 18),
 658 => to_signed(0, 18),
 659 => to_signed(0, 18),
 660 => to_signed(0, 18),
 661 => to_signed(0, 18),
 662 => to_signed(0, 18),
 663 => to_signed(0, 18),
 664 => to_signed(0, 18),
 665 => to_signed(0, 18),
 666 => to_signed(0, 18),
 667 => to_signed(0, 18),
 668 => to_signed(0, 18),
 669 => to_signed(0, 18),
 670 => to_signed(0, 18),
 671 => to_signed(0, 18),
 672 => to_signed(0, 18),
 673 => to_signed(0, 18),
 674 => to_signed(0, 18),
 675 => to_signed(0, 18),
 676 => to_signed(0, 18),
 677 => to_signed(0, 18),
 678 => to_signed(0, 18),
 679 => to_signed(0, 18),
 680 => to_signed(0, 18),
 681 => to_signed(0, 18),
 682 => to_signed(0, 18),
 683 => to_signed(0, 18),
 684 => to_signed(0, 18),
 685 => to_signed(0, 18),
 686 => to_signed(0, 18),
 687 => to_signed(0, 18),
 688 => to_signed(0, 18),
 689 => to_signed(0, 18),
 690 => to_signed(0, 18),
 691 => to_signed(0, 18),
 692 => to_signed(0, 18),
 693 => to_signed(0, 18),
 694 => to_signed(0, 18),
 695 => to_signed(0, 18),
 696 => to_signed(0, 18),
 697 => to_signed(0, 18),
 698 => to_signed(0, 18),
 699 => to_signed(0, 18),
 700 => to_signed(0, 18),
 701 => to_signed(0, 18),
 702 => to_signed(0, 18),
 703 => to_signed(0, 18),
 704 => to_signed(0, 18),
 705 => to_signed(0, 18),
 706 => to_signed(0, 18),
 707 => to_signed(0, 18),
 708 => to_signed(0, 18),
 709 => to_signed(0, 18),
 710 => to_signed(0, 18),
 711 => to_signed(0, 18),
 712 => to_signed(0, 18),
 713 => to_signed(0, 18),
 714 => to_signed(0, 18),
 715 => to_signed(0, 18),
 716 => to_signed(0, 18),
 717 => to_signed(0, 18),
 718 => to_signed(0, 18),
 719 => to_signed(0, 18),
 720 => to_signed(0, 18),
 721 => to_signed(0, 18),
 722 => to_signed(0, 18),
 723 => to_signed(0, 18),
 724 => to_signed(0, 18),
 725 => to_signed(0, 18),
 726 => to_signed(0, 18),
 727 => to_signed(0, 18),
 728 => to_signed(0, 18),
 729 => to_signed(0, 18),
 730 => to_signed(0, 18),
 731 => to_signed(0, 18),
 732 => to_signed(0, 18),
 733 => to_signed(0, 18),
 734 => to_signed(0, 18),
 735 => to_signed(0, 18),
 736 => to_signed(0, 18),
 737 => to_signed(0, 18),
 738 => to_signed(0, 18),
 739 => to_signed(0, 18),
 740 => to_signed(0, 18),
 741 => to_signed(0, 18),
 742 => to_signed(0, 18),
 743 => to_signed(0, 18),
 744 => to_signed(0, 18),
 745 => to_signed(0, 18),
 746 => to_signed(0, 18),
 747 => to_signed(0, 18),
 748 => to_signed(0, 18),
 749 => to_signed(0, 18),
 750 => to_signed(0, 18),
 751 => to_signed(0, 18),
 752 => to_signed(0, 18),
 753 => to_signed(0, 18),
 754 => to_signed(0, 18),
 755 => to_signed(0, 18),
 756 => to_signed(0, 18),
 757 => to_signed(0, 18),
 758 => to_signed(0, 18),
 759 => to_signed(0, 18),
 760 => to_signed(0, 18),
 761 => to_signed(0, 18),
 762 => to_signed(0, 18),
 763 => to_signed(0, 18),
 764 => to_signed(0, 18),
 765 => to_signed(0, 18),
 766 => to_signed(0, 18),
 767 => to_signed(0, 18),
 768 => to_signed(0, 18),
 769 => to_signed(0, 18),
 770 => to_signed(0, 18),
 771 => to_signed(0, 18),
 772 => to_signed(0, 18),
 773 => to_signed(0, 18),
 774 => to_signed(0, 18),
 775 => to_signed(0, 18),
 776 => to_signed(0, 18),
 777 => to_signed(0, 18),
 778 => to_signed(0, 18),
 779 => to_signed(0, 18),
 780 => to_signed(0, 18),
 781 => to_signed(0, 18),
 782 => to_signed(0, 18),
 783 => to_signed(0, 18),
 784 => to_signed(0, 18),
 785 => to_signed(0, 18),
 786 => to_signed(0, 18),
 787 => to_signed(0, 18),
 788 => to_signed(0, 18),
 789 => to_signed(0, 18),
 790 => to_signed(0, 18),
 791 => to_signed(0, 18),
 792 => to_signed(0, 18),
 793 => to_signed(0, 18),
 794 => to_signed(0, 18),
 795 => to_signed(0, 18),
 796 => to_signed(0, 18),
 797 => to_signed(0, 18),
 798 => to_signed(0, 18),
 799 => to_signed(0, 18),
 800 => to_signed(0, 18),
 801 => to_signed(0, 18),
 802 => to_signed(0, 18),
 803 => to_signed(0, 18),
 804 => to_signed(0, 18),
 805 => to_signed(0, 18),
 806 => to_signed(0, 18),
 807 => to_signed(0, 18),
 808 => to_signed(0, 18),
 809 => to_signed(0, 18),
 810 => to_signed(0, 18),
 811 => to_signed(0, 18),
 812 => to_signed(0, 18),
 813 => to_signed(0, 18),
 814 => to_signed(0, 18),
 815 => to_signed(0, 18),
 816 => to_signed(0, 18),
 817 => to_signed(0, 18),
 818 => to_signed(0, 18),
 819 => to_signed(0, 18),
 820 => to_signed(0, 18),
 821 => to_signed(0, 18),
 822 => to_signed(0, 18),
 823 => to_signed(0, 18),
 824 => to_signed(0, 18),
 825 => to_signed(0, 18),
 826 => to_signed(0, 18),
 827 => to_signed(0, 18),
 828 => to_signed(0, 18),
 829 => to_signed(0, 18),
 830 => to_signed(0, 18),
 831 => to_signed(0, 18),
 832 => to_signed(0, 18),
 833 => to_signed(0, 18),
 834 => to_signed(0, 18),
 835 => to_signed(0, 18),
 836 => to_signed(0, 18),
 837 => to_signed(0, 18),
 838 => to_signed(0, 18),
 839 => to_signed(0, 18),
 840 => to_signed(0, 18),
 841 => to_signed(0, 18),
 842 => to_signed(0, 18),
 843 => to_signed(0, 18),
 844 => to_signed(0, 18),
 845 => to_signed(0, 18),
 846 => to_signed(0, 18),
 847 => to_signed(0, 18),
 848 => to_signed(0, 18),
 849 => to_signed(0, 18),
 850 => to_signed(0, 18),
 851 => to_signed(0, 18),
 852 => to_signed(0, 18),
 853 => to_signed(0, 18),
 854 => to_signed(0, 18),
 855 => to_signed(0, 18),
 856 => to_signed(0, 18),
 857 => to_signed(0, 18),
 858 => to_signed(0, 18),
 859 => to_signed(0, 18),
 860 => to_signed(0, 18),
 861 => to_signed(0, 18),
 862 => to_signed(0, 18),
 863 => to_signed(0, 18),
 864 => to_signed(0, 18),
 865 => to_signed(0, 18),
 866 => to_signed(0, 18),
 867 => to_signed(0, 18),
 868 => to_signed(0, 18),
 869 => to_signed(0, 18),
 870 => to_signed(0, 18),
 871 => to_signed(0, 18),
 872 => to_signed(0, 18),
 873 => to_signed(0, 18),
 874 => to_signed(0, 18),
 875 => to_signed(0, 18),
 876 => to_signed(0, 18),
 877 => to_signed(0, 18),
 878 => to_signed(0, 18),
 879 => to_signed(0, 18),
 880 => to_signed(0, 18),
 881 => to_signed(0, 18),
 882 => to_signed(0, 18),
 883 => to_signed(0, 18),
 884 => to_signed(0, 18),
 885 => to_signed(0, 18),
 886 => to_signed(0, 18),
 887 => to_signed(0, 18),
 888 => to_signed(0, 18),
 889 => to_signed(0, 18),
 890 => to_signed(0, 18),
 891 => to_signed(0, 18),
 892 => to_signed(0, 18),
 893 => to_signed(0, 18),
 894 => to_signed(0, 18),
 895 => to_signed(0, 18),
 896 => to_signed(0, 18),
 897 => to_signed(0, 18),
 898 => to_signed(0, 18),
 899 => to_signed(0, 18));

begin

DUT : test_iir
port map (
	CLK => CLK,
	DATA_IN => DATA_IN,
	DATA_IN_VAL => DATA_IN_VAL,
	SRST => SRST,
	DATA_OUT => DATA_OUT,
	DATA_OUT_VAL => DATA_OUT_VAL
	);

CLK <= not CLK after CLK_PERIOD/2;

STIMULUS_DATA_IN_PROCESS : process
procedure tic (nb_cycles : natural := 1) is
begin
	for I in 1 to nb_cycles loop
		wait until rising_edge(CLK);
	end loop;
end procedure;

begin
	DATA_IN_VAL <= '0';
	DATA_IN <= to_signed(0, DATA_IN'length);
	tic;
	SRST <= '1';
	tic;
	SRST <= '0';
	tic;
	assert DATA_OUT = 0 report "DATA_OUT must be 0 after a reset";
	assert DATA_OUT_VAL = '0' report "DATA_OUT_VAL must be 0 after a reset";
	tic;
	for I in DATA_IN_ARRAY'range loop
		DATA_IN_VAL <= '1';
		DATA_IN <= DATA_IN_ARRAY(I);
		tic;
	end loop;
	DATA_IN_VAL <= '0';
	tic(20); -- Make sure all data has been processed
	SRST <= '1';
	tic;
	SRST <= '0';
	tic;
	assert DATA_OUT = 0 report "DATA_OUT must be 0 after a reset";
	assert DATA_OUT_VAL = '0' report "DATA_OUT_VAL must be 0 after a reset";
	tic;	
	for I in DATA_IN_ARRAY'range loop
		DATA_IN_VAL <= '1';
		DATA_IN <= DATA_IN_ARRAY(I);
		tic;
		DATA_IN_VAL <= '0'; -- Now we simulate, new data on every other clock cycle
		tic;
	end loop;
	tic(20);
	std.env.finish;
end process;

STIMULUS_DATA_OUT_PROCESS : process
variable cnt : natural := 0;
procedure tic (nb_cycles : natural := 1) is
begin
	for I in 1 to nb_cycles loop
		wait until rising_edge(CLK);
	end loop;
end procedure;

begin
	wait until rising_edge(CLK);
	if (DATA_OUT_VAL = '1') then
		assert (DATA_OUT = DATA_OUT_ARRAY(cnt)) report "Error data out = " & integer'image(to_integer(DATA_OUT)) & "Should be " & integer'image(to_integer(DATA_OUT_ARRAY(cnt))) & " on sample " & integer'image(cnt) severity error;
		cnt := cnt + 1;
	elsif (SRST = '1') then
		cnt := 0;
	end if;
			
	
	
end process;

	
end architecture TB;

